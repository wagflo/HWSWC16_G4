-- raytracing.vhd

-- Generated using ACDS version 16.0 222

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity raytracing is
	port (
		altpll_0_areset_conduit_export : in    std_logic                     := '0';             -- altpll_0_areset_conduit.export
		altpll_0_locked_conduit_export : out   std_logic;                                        -- altpll_0_locked_conduit.export
		altpll_c4_conduit_export       : out   std_logic;                                        --       altpll_c4_conduit.export
		clk_clk                        : in    std_logic                     := '0';             --                     clk.clk
		ltm_vid_data                   : out   std_logic_vector(23 downto 0);                    --                     ltm.vid_data
		ltm_underflow                  : out   std_logic;                                        --                        .underflow
		ltm_vid_datavalid              : out   std_logic;                                        --                        .vid_datavalid
		ltm_vid_v_sync                 : out   std_logic;                                        --                        .vid_v_sync
		ltm_vid_h_sync                 : out   std_logic;                                        --                        .vid_h_sync
		ltm_vid_f                      : out   std_logic;                                        --                        .vid_f
		ltm_vid_h                      : out   std_logic;                                        --                        .vid_h
		ltm_vid_v                      : out   std_logic;                                        --                        .vid_v
		ltm_clk_clk                    : out   std_logic;                                        --                 ltm_clk.clk
		reset_reset_n                  : in    std_logic                     := '0';             --                   reset.reset_n
		sdram_addr                     : out   std_logic_vector(12 downto 0);                    --                   sdram.addr
		sdram_ba                       : out   std_logic_vector(1 downto 0);                     --                        .ba
		sdram_cas_n                    : out   std_logic;                                        --                        .cas_n
		sdram_cke                      : out   std_logic;                                        --                        .cke
		sdram_cs_n                     : out   std_logic;                                        --                        .cs_n
		sdram_dq                       : inout std_logic_vector(31 downto 0) := (others => '0'); --                        .dq
		sdram_dqm                      : out   std_logic_vector(3 downto 0);                     --                        .dqm
		sdram_ras_n                    : out   std_logic;                                        --                        .ras_n
		sdram_we_n                     : out   std_logic;                                        --                        .we_n
		sdram_clk_clk                  : out   std_logic                                         --               sdram_clk.clk
	);
end entity raytracing;

architecture rtl of raytracing is
	component raytracing_altpll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			c4                 : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component raytracing_altpll;

	component alt_vipvfr131_vfr is
		generic (
			BITS_PER_PIXEL_PER_COLOR_PLANE : integer := 8;
			NUMBER_OF_CHANNELS_IN_PARALLEL : integer := 3;
			NUMBER_OF_CHANNELS_IN_SEQUENCE : integer := 1;
			MAX_IMAGE_WIDTH                : integer := 640;
			MAX_IMAGE_HEIGHT               : integer := 480;
			MEM_PORT_WIDTH                 : integer := 256;
			RMASTER_FIFO_DEPTH             : integer := 64;
			RMASTER_BURST_TARGET           : integer := 32;
			CLOCKS_ARE_SEPARATE            : integer := 1
		);
		port (
			clock                : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_clock         : in  std_logic                     := 'X';             -- clk
			master_reset         : in  std_logic                     := 'X';             -- reset
			slave_address        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			slave_irq            : out std_logic;                                        -- irq
			dout_data            : out std_logic_vector(23 downto 0);                    -- data
			dout_valid           : out std_logic;                                        -- valid
			dout_ready           : in  std_logic                     := 'X';             -- ready
			dout_startofpacket   : out std_logic;                                        -- startofpacket
			dout_endofpacket     : out std_logic;                                        -- endofpacket
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_burstcount    : out std_logic_vector(5 downto 0);                     -- burstcount
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X'              -- waitrequest
		);
	end component alt_vipvfr131_vfr;

	component raytracing_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component raytracing_jtag_uart;

	component alt_vipitc131_IS2Vid is
		generic (
			NUMBER_OF_COLOUR_PLANES       : integer := 3;
			COLOUR_PLANES_ARE_IN_PARALLEL : integer := 1;
			BPS                           : integer := 8;
			INTERLACED                    : integer := 0;
			H_ACTIVE_PIXELS               : integer := 1920;
			V_ACTIVE_LINES                : integer := 1200;
			ACCEPT_COLOURS_IN_SEQ         : integer := 0;
			FIFO_DEPTH                    : integer := 1920;
			CLOCKS_ARE_SAME               : integer := 0;
			USE_CONTROL                   : integer := 0;
			NO_OF_MODES                   : integer := 1;
			THRESHOLD                     : integer := 1919;
			STD_WIDTH                     : integer := 1;
			GENERATE_SYNC                 : integer := 0;
			USE_EMBEDDED_SYNCS            : integer := 0;
			AP_LINE                       : integer := 0;
			V_BLANK                       : integer := 0;
			H_BLANK                       : integer := 0;
			H_SYNC_LENGTH                 : integer := 44;
			H_FRONT_PORCH                 : integer := 88;
			H_BACK_PORCH                  : integer := 148;
			V_SYNC_LENGTH                 : integer := 5;
			V_FRONT_PORCH                 : integer := 4;
			V_BACK_PORCH                  : integer := 36;
			F_RISING_EDGE                 : integer := 0;
			F_FALLING_EDGE                : integer := 0;
			FIELD0_V_RISING_EDGE          : integer := 0;
			FIELD0_V_BLANK                : integer := 0;
			FIELD0_V_SYNC_LENGTH          : integer := 0;
			FIELD0_V_FRONT_PORCH          : integer := 0;
			FIELD0_V_BACK_PORCH           : integer := 0;
			ANC_LINE                      : integer := 0;
			FIELD0_ANC_LINE               : integer := 0
		);
		port (
			is_clk        : in  std_logic                     := 'X';             -- clk
			rst           : in  std_logic                     := 'X';             -- reset
			is_data       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			is_valid      : in  std_logic                     := 'X';             -- valid
			is_ready      : out std_logic;                                        -- ready
			is_sop        : in  std_logic                     := 'X';             -- startofpacket
			is_eop        : in  std_logic                     := 'X';             -- endofpacket
			vid_data      : out std_logic_vector(23 downto 0);                    -- export
			underflow     : out std_logic;                                        -- export
			vid_datavalid : out std_logic;                                        -- export
			vid_v_sync    : out std_logic;                                        -- export
			vid_h_sync    : out std_logic;                                        -- export
			vid_f         : out std_logic;                                        -- export
			vid_h         : out std_logic;                                        -- export
			vid_v         : out std_logic                                         -- export
		);
	end component alt_vipitc131_IS2Vid;

	component raytracing_mm is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			res_n            : in  std_logic                     := 'X';             -- reset
			address          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			write            : in  std_logic                     := 'X';             -- write
			writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			master_address   : out std_logic_vector(31 downto 0);                    -- address
			master_write     : out std_logic;                                        -- write
			master_colordata : out std_logic_vector(31 downto 0);                    -- writedata
			slave_waitreq    : in  std_logic                     := 'X'              -- waitrequest
		);
	end component raytracing_mm;

	component raytracing_nios2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component raytracing_nios2;

	component raytracing_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component raytracing_onchip_ram;

	component raytracing_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component raytracing_sdram;

	component raytracing_systimer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component raytracing_systimer;

	component raytracing_mm_interconnect_0 is
		port (
			altpll_c0_clk                                              : in  std_logic                     := 'X';             -- clk
			altpll_c1_clk                                              : in  std_logic                     := 'X';             -- clk
			altpll_c3_clk                                              : in  std_logic                     := 'X';             -- clk
			clk_50_clk_clk                                             : in  std_logic                     := 'X';             -- clk
			altpll_inclk_interface_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			framereader_clock_master_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			framereader_clock_reset_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			mm_raytracing_0_reset_sink_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			nios2_reset_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			framereader_avalon_master_address                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			framereader_avalon_master_waitrequest                      : out std_logic;                                        -- waitrequest
			framereader_avalon_master_burstcount                       : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- burstcount
			framereader_avalon_master_read                             : in  std_logic                     := 'X';             -- read
			framereader_avalon_master_readdata                         : out std_logic_vector(31 downto 0);                    -- readdata
			framereader_avalon_master_readdatavalid                    : out std_logic;                                        -- readdatavalid
			mm_raytracing_0_mm_sdram_master_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			mm_raytracing_0_mm_sdram_master_waitrequest                : out std_logic;                                        -- waitrequest
			mm_raytracing_0_mm_sdram_master_write                      : in  std_logic                     := 'X';             -- write
			mm_raytracing_0_mm_sdram_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_address                                  : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_data_master_waitrequest                              : out std_logic;                                        -- waitrequest
			nios2_data_master_byteenable                               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_data_master_read                                     : in  std_logic                     := 'X';             -- read
			nios2_data_master_readdata                                 : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_data_master_readdatavalid                            : out std_logic;                                        -- readdatavalid
			nios2_data_master_write                                    : in  std_logic                     := 'X';             -- write
			nios2_data_master_writedata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_debugaccess                              : in  std_logic                     := 'X';             -- debugaccess
			nios2_instruction_master_address                           : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_instruction_master_waitrequest                       : out std_logic;                                        -- waitrequest
			nios2_instruction_master_read                              : in  std_logic                     := 'X';             -- read
			nios2_instruction_master_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_instruction_master_readdatavalid                     : out std_logic;                                        -- readdatavalid
			altpll_pll_slave_address                                   : out std_logic_vector(1 downto 0);                     -- address
			altpll_pll_slave_write                                     : out std_logic;                                        -- write
			altpll_pll_slave_read                                      : out std_logic;                                        -- read
			altpll_pll_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_pll_slave_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			framereader_avalon_slave_address                           : out std_logic_vector(4 downto 0);                     -- address
			framereader_avalon_slave_write                             : out std_logic;                                        -- write
			framereader_avalon_slave_read                              : out std_logic;                                        -- read
			framereader_avalon_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			framereader_avalon_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                          : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                           : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                     : out std_logic;                                        -- chipselect
			mm_raytracing_0_mm_nios_slave_address                      : out std_logic_vector(15 downto 0);                    -- address
			mm_raytracing_0_mm_nios_slave_write                        : out std_logic;                                        -- write
			mm_raytracing_0_mm_nios_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_debug_mem_slave_address                              : out std_logic_vector(8 downto 0);                     -- address
			nios2_debug_mem_slave_write                                : out std_logic;                                        -- write
			nios2_debug_mem_slave_read                                 : out std_logic;                                        -- read
			nios2_debug_mem_slave_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_debug_mem_slave_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_debug_mem_slave_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_debug_mem_slave_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			nios2_debug_mem_slave_debugaccess                          : out std_logic;                                        -- debugaccess
			onchip_ram_s1_address                                      : out std_logic_vector(15 downto 0);                    -- address
			onchip_ram_s1_write                                        : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                                   : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                        : out std_logic;                                        -- clken
			sdram_s1_address                                           : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                             : out std_logic;                                        -- write
			sdram_s1_read                                              : out std_logic;                                        -- read
			sdram_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_s1_byteenable                                        : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                     : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                       : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                        : out std_logic;                                        -- chipselect
			systimer_s1_address                                        : out std_logic_vector(3 downto 0);                     -- address
			systimer_s1_write                                          : out std_logic;                                        -- write
			systimer_s1_readdata                                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			systimer_s1_writedata                                      : out std_logic_vector(15 downto 0);                    -- writedata
			systimer_s1_chipselect                                     : out std_logic                                         -- chipselect
		);
	end component raytracing_mm_interconnect_0;

	component raytracing_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component raytracing_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component raytracing_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component raytracing_rst_controller;

	component raytracing_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component raytracing_rst_controller_002;

	component raytracing_rst_controller_004 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component raytracing_rst_controller_004;

	signal framereader_avalon_streaming_source_valid                     : std_logic;                     -- framereader:dout_valid -> ltm:is_valid
	signal framereader_avalon_streaming_source_data                      : std_logic_vector(23 downto 0); -- framereader:dout_data -> ltm:is_data
	signal framereader_avalon_streaming_source_ready                     : std_logic;                     -- ltm:is_ready -> framereader:dout_ready
	signal framereader_avalon_streaming_source_startofpacket             : std_logic;                     -- framereader:dout_startofpacket -> ltm:is_sop
	signal framereader_avalon_streaming_source_endofpacket               : std_logic;                     -- framereader:dout_endofpacket -> ltm:is_eop
	signal altpll_c0_clk                                                 : std_logic;                     -- altpll:c0 -> [framereader:master_clock, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, mm_interconnect_0:altpll_c0_clk, nios2:clk, onchip_ram:clk, rst_controller_002:clk, rst_controller_004:clk, sdram:clk, systimer:clk]
	signal altpll_c1_clk                                                 : std_logic;                     -- altpll:c1 -> [ltm_clk_clk, framereader:clock, irq_synchronizer:receiver_clk, ltm:is_clk, mm_interconnect_0:altpll_c1_clk, rst_controller_001:clk]
	signal altpll_c3_clk                                                 : std_logic;                     -- altpll:c3 -> [mm_interconnect_0:altpll_c3_clk, mm_raytracing_0:clk, rst_controller_003:clk]
	signal framereader_avalon_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:framereader_avalon_master_readdata -> framereader:master_readdata
	signal framereader_avalon_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:framereader_avalon_master_waitrequest -> framereader:master_waitrequest
	signal framereader_avalon_master_address                             : std_logic_vector(31 downto 0); -- framereader:master_address -> mm_interconnect_0:framereader_avalon_master_address
	signal framereader_avalon_master_read                                : std_logic;                     -- framereader:master_read -> mm_interconnect_0:framereader_avalon_master_read
	signal framereader_avalon_master_readdatavalid                       : std_logic;                     -- mm_interconnect_0:framereader_avalon_master_readdatavalid -> framereader:master_readdatavalid
	signal framereader_avalon_master_burstcount                          : std_logic_vector(5 downto 0);  -- framereader:master_burstcount -> mm_interconnect_0:framereader_avalon_master_burstcount
	signal nios2_data_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	signal nios2_data_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	signal nios2_data_master_debugaccess                                 : std_logic;                     -- nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	signal nios2_data_master_address                                     : std_logic_vector(27 downto 0); -- nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	signal nios2_data_master_byteenable                                  : std_logic_vector(3 downto 0);  -- nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	signal nios2_data_master_read                                        : std_logic;                     -- nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	signal nios2_data_master_readdatavalid                               : std_logic;                     -- mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	signal nios2_data_master_write                                       : std_logic;                     -- nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	signal nios2_data_master_writedata                                   : std_logic_vector(31 downto 0); -- nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	signal mm_raytracing_0_mm_sdram_master_waitrequest                   : std_logic;                     -- mm_interconnect_0:mm_raytracing_0_mm_sdram_master_waitrequest -> mm_raytracing_0:slave_waitreq
	signal mm_raytracing_0_mm_sdram_master_address                       : std_logic_vector(31 downto 0); -- mm_raytracing_0:master_address -> mm_interconnect_0:mm_raytracing_0_mm_sdram_master_address
	signal mm_raytracing_0_mm_sdram_master_write                         : std_logic;                     -- mm_raytracing_0:master_write -> mm_interconnect_0:mm_raytracing_0_mm_sdram_master_write
	signal mm_raytracing_0_mm_sdram_master_writedata                     : std_logic_vector(31 downto 0); -- mm_raytracing_0:master_colordata -> mm_interconnect_0:mm_raytracing_0_mm_sdram_master_writedata
	signal nios2_instruction_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	signal nios2_instruction_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	signal nios2_instruction_master_address                              : std_logic_vector(26 downto 0); -- nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	signal nios2_instruction_master_read                                 : std_logic;                     -- nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	signal nios2_instruction_master_readdatavalid                        : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	signal mm_interconnect_0_sdram_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                           : std_logic_vector(31 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                        : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                            : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                               : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                      : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                              : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_framereader_avalon_slave_readdata           : std_logic_vector(31 downto 0); -- framereader:slave_readdata -> mm_interconnect_0:framereader_avalon_slave_readdata
	signal mm_interconnect_0_framereader_avalon_slave_address            : std_logic_vector(4 downto 0);  -- mm_interconnect_0:framereader_avalon_slave_address -> framereader:slave_address
	signal mm_interconnect_0_framereader_avalon_slave_read               : std_logic;                     -- mm_interconnect_0:framereader_avalon_slave_read -> framereader:slave_read
	signal mm_interconnect_0_framereader_avalon_slave_write              : std_logic;                     -- mm_interconnect_0:framereader_avalon_slave_write -> framereader:slave_write
	signal mm_interconnect_0_framereader_avalon_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:framereader_avalon_slave_writedata -> framereader:slave_writedata
	signal mm_interconnect_0_nios2_debug_mem_slave_readdata              : std_logic_vector(31 downto 0); -- nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_debug_mem_slave_waitrequest           : std_logic;                     -- nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_debug_mem_slave_debugaccess           : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_debug_mem_slave_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	signal mm_interconnect_0_nios2_debug_mem_slave_read                  : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	signal mm_interconnect_0_nios2_debug_mem_slave_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_debug_mem_slave_write                 : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	signal mm_interconnect_0_nios2_debug_mem_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	signal mm_interconnect_0_mm_raytracing_0_mm_nios_slave_address       : std_logic_vector(15 downto 0); -- mm_interconnect_0:mm_raytracing_0_mm_nios_slave_address -> mm_raytracing_0:address
	signal mm_interconnect_0_mm_raytracing_0_mm_nios_slave_write         : std_logic;                     -- mm_interconnect_0:mm_raytracing_0_mm_nios_slave_write -> mm_raytracing_0:write
	signal mm_interconnect_0_mm_raytracing_0_mm_nios_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_raytracing_0_mm_nios_slave_writedata -> mm_raytracing_0:writedata
	signal mm_interconnect_0_altpll_pll_slave_readdata                   : std_logic_vector(31 downto 0); -- altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	signal mm_interconnect_0_altpll_pll_slave_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	signal mm_interconnect_0_altpll_pll_slave_read                       : std_logic;                     -- mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	signal mm_interconnect_0_altpll_pll_slave_write                      : std_logic;                     -- mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	signal mm_interconnect_0_altpll_pll_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	signal mm_interconnect_0_systimer_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:systimer_s1_chipselect -> systimer:chipselect
	signal mm_interconnect_0_systimer_s1_readdata                        : std_logic_vector(15 downto 0); -- systimer:readdata -> mm_interconnect_0:systimer_s1_readdata
	signal mm_interconnect_0_systimer_s1_address                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:systimer_s1_address -> systimer:address
	signal mm_interconnect_0_systimer_s1_write                           : std_logic;                     -- mm_interconnect_0:systimer_s1_write -> mm_interconnect_0_systimer_s1_write:in
	signal mm_interconnect_0_systimer_s1_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:systimer_s1_writedata -> systimer:writedata
	signal mm_interconnect_0_onchip_ram_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- systimer:irq -> irq_mapper:receiver2_irq
	signal nios2_irq_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2:irq
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                 : std_logic_vector(0 downto 0);  -- framereader:slave_irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [framereader:reset, irq_synchronizer:receiver_reset, ltm:rst, mm_interconnect_0:framereader_clock_reset_reset_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [framereader:master_reset, mm_interconnect_0:framereader_clock_master_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_002_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_002_reset_out_reset_req                        : std_logic;                     -- rst_controller_002:reset_req -> [onchip_ram:reset_req, rst_translator:reset_req_in]
	signal rst_controller_003_reset_out_reset                            : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:mm_raytracing_0_reset_sink_reset_bridge_in_reset_reset, mm_raytracing_0:res_n]
	signal rst_controller_004_reset_out_reset                            : std_logic;                     -- rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, rst_controller_004_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_004_reset_out_reset_req                        : std_logic;                     -- rst_controller_004:reset_req -> [nios2:reset_req, rst_translator_001:reset_req_in]
	signal nios2_debug_reset_request_reset                               : std_logic;                     -- nios2:debug_reset_request -> rst_controller_004:reset_in1
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0]
	signal mm_interconnect_0_sdram_s1_read_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv               : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_systimer_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_systimer_s1_write:inv -> systimer:write_n
	signal rst_controller_002_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [jtag_uart:rst_n, sdram:reset_n, systimer:reset_n]
	signal rst_controller_004_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_004_reset_out_reset:inv -> nios2:reset_n

begin

	altpll : component raytracing_altpll
		port map (
			clk                => clk_clk,                                      --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,               -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_pll_slave_writedata, --                      .writedata
			c0                 => altpll_c0_clk,                                --                    c0.clk
			c1                 => altpll_c1_clk,                                --                    c1.clk
			c2                 => sdram_clk_clk,                                --                    c2.clk
			c3                 => altpll_c3_clk,                                --                    c3.clk
			areset             => altpll_0_areset_conduit_export,               --        areset_conduit.export
			locked             => altpll_0_locked_conduit_export,               --        locked_conduit.export
			c4                 => altpll_c4_conduit_export,                     --            c4_conduit.export
			scandone           => open,                                         --           (terminated)
			scandataout        => open,                                         --           (terminated)
			phasedone          => open,                                         --           (terminated)
			phasecounterselect => "0000",                                       --           (terminated)
			phaseupdown        => '0',                                          --           (terminated)
			phasestep          => '0',                                          --           (terminated)
			scanclk            => '0',                                          --           (terminated)
			scanclkena         => '0',                                          --           (terminated)
			scandata           => '0',                                          --           (terminated)
			configupdate       => '0'                                           --           (terminated)
		);

	framereader : component alt_vipvfr131_vfr
		generic map (
			BITS_PER_PIXEL_PER_COLOR_PLANE => 8,
			NUMBER_OF_CHANNELS_IN_PARALLEL => 3,
			NUMBER_OF_CHANNELS_IN_SEQUENCE => 1,
			MAX_IMAGE_WIDTH                => 800,
			MAX_IMAGE_HEIGHT               => 480,
			MEM_PORT_WIDTH                 => 32,
			RMASTER_FIFO_DEPTH             => 64,
			RMASTER_BURST_TARGET           => 32,
			CLOCKS_ARE_SEPARATE            => 1
		)
		port map (
			clock                => altpll_c1_clk,                                        --             clock_reset.clk
			reset                => rst_controller_001_reset_out_reset,                   --       clock_reset_reset.reset
			master_clock         => altpll_c0_clk,                                        --            clock_master.clk
			master_reset         => rst_controller_002_reset_out_reset,                   --      clock_master_reset.reset
			slave_address        => mm_interconnect_0_framereader_avalon_slave_address,   --            avalon_slave.address
			slave_write          => mm_interconnect_0_framereader_avalon_slave_write,     --                        .write
			slave_writedata      => mm_interconnect_0_framereader_avalon_slave_writedata, --                        .writedata
			slave_read           => mm_interconnect_0_framereader_avalon_slave_read,      --                        .read
			slave_readdata       => mm_interconnect_0_framereader_avalon_slave_readdata,  --                        .readdata
			slave_irq            => irq_synchronizer_receiver_irq(0),                     --        interrupt_sender.irq
			dout_data            => framereader_avalon_streaming_source_data,             -- avalon_streaming_source.data
			dout_valid           => framereader_avalon_streaming_source_valid,            --                        .valid
			dout_ready           => framereader_avalon_streaming_source_ready,            --                        .ready
			dout_startofpacket   => framereader_avalon_streaming_source_startofpacket,    --                        .startofpacket
			dout_endofpacket     => framereader_avalon_streaming_source_endofpacket,      --                        .endofpacket
			master_address       => framereader_avalon_master_address,                    --           avalon_master.address
			master_burstcount    => framereader_avalon_master_burstcount,                 --                        .burstcount
			master_readdata      => framereader_avalon_master_readdata,                   --                        .readdata
			master_read          => framereader_avalon_master_read,                       --                        .read
			master_readdatavalid => framereader_avalon_master_readdatavalid,              --                        .readdatavalid
			master_waitrequest   => framereader_avalon_master_waitrequest                 --                        .waitrequest
		);

	jtag_uart : component raytracing_jtag_uart
		port map (
			clk            => altpll_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	ltm : component alt_vipitc131_IS2Vid
		generic map (
			NUMBER_OF_COLOUR_PLANES       => 3,
			COLOUR_PLANES_ARE_IN_PARALLEL => 1,
			BPS                           => 8,
			INTERLACED                    => 0,
			H_ACTIVE_PIXELS               => 800,
			V_ACTIVE_LINES                => 480,
			ACCEPT_COLOURS_IN_SEQ         => 0,
			FIFO_DEPTH                    => 1024,
			CLOCKS_ARE_SAME               => 1,
			USE_CONTROL                   => 0,
			NO_OF_MODES                   => 1,
			THRESHOLD                     => 1023,
			STD_WIDTH                     => 1,
			GENERATE_SYNC                 => 0,
			USE_EMBEDDED_SYNCS            => 0,
			AP_LINE                       => 0,
			V_BLANK                       => 0,
			H_BLANK                       => 0,
			H_SYNC_LENGTH                 => 1,
			H_FRONT_PORCH                 => 40,
			H_BACK_PORCH                  => 216,
			V_SYNC_LENGTH                 => 1,
			V_FRONT_PORCH                 => 10,
			V_BACK_PORCH                  => 35,
			F_RISING_EDGE                 => 0,
			F_FALLING_EDGE                => 0,
			FIELD0_V_RISING_EDGE          => 0,
			FIELD0_V_BLANK                => 0,
			FIELD0_V_SYNC_LENGTH          => 0,
			FIELD0_V_FRONT_PORCH          => 0,
			FIELD0_V_BACK_PORCH           => 0,
			ANC_LINE                      => 0,
			FIELD0_ANC_LINE               => 0
		)
		port map (
			is_clk        => altpll_c1_clk,                                     --       is_clk_rst.clk
			rst           => rst_controller_001_reset_out_reset,                -- is_clk_rst_reset.reset
			is_data       => framereader_avalon_streaming_source_data,          --              din.data
			is_valid      => framereader_avalon_streaming_source_valid,         --                 .valid
			is_ready      => framereader_avalon_streaming_source_ready,         --                 .ready
			is_sop        => framereader_avalon_streaming_source_startofpacket, --                 .startofpacket
			is_eop        => framereader_avalon_streaming_source_endofpacket,   --                 .endofpacket
			vid_data      => ltm_vid_data,                                      --    clocked_video.export
			underflow     => ltm_underflow,                                     --                 .export
			vid_datavalid => ltm_vid_datavalid,                                 --                 .export
			vid_v_sync    => ltm_vid_v_sync,                                    --                 .export
			vid_h_sync    => ltm_vid_h_sync,                                    --                 .export
			vid_f         => ltm_vid_f,                                         --                 .export
			vid_h         => ltm_vid_h,                                         --                 .export
			vid_v         => ltm_vid_v                                          --                 .export
		);

	mm_raytracing_0 : component raytracing_mm
		port map (
			clk              => altpll_c3_clk,                                             --      clock_sink.clk
			res_n            => rst_controller_003_reset_out_reset,                        --      reset_sink.reset
			address          => mm_interconnect_0_mm_raytracing_0_mm_nios_slave_address,   --   mm_nios_slave.address
			write            => mm_interconnect_0_mm_raytracing_0_mm_nios_slave_write,     --                .write
			writedata        => mm_interconnect_0_mm_raytracing_0_mm_nios_slave_writedata, --                .writedata
			master_address   => mm_raytracing_0_mm_sdram_master_address,                   -- mm_sdram_master.address
			master_write     => mm_raytracing_0_mm_sdram_master_write,                     --                .write
			master_colordata => mm_raytracing_0_mm_sdram_master_writedata,                 --                .writedata
			slave_waitreq    => mm_raytracing_0_mm_sdram_master_waitrequest                --                .waitrequest
		);

	nios2 : component raytracing_nios2
		port map (
			clk                                 => altpll_c0_clk,                                       --                       clk.clk
			reset_n                             => rst_controller_004_reset_out_reset_ports_inv,        --                     reset.reset_n
			reset_req                           => rst_controller_004_reset_out_reset_req,              --                          .reset_req
			d_address                           => nios2_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_data_master_read,                              --                          .read
			d_readdata                          => nios2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_data_master_write,                             --                          .write
			d_writedata                         => nios2_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	onchip_ram : component raytracing_onchip_ram
		port map (
			clk        => altpll_c0_clk,                              --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_002_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_002_reset_out_reset_req      --       .reset_req
		);

	sdram : component raytracing_sdram
		port map (
			clk            => altpll_c0_clk,                                   --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,    -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	systimer : component raytracing_systimer
		port map (
			clk        => altpll_c0_clk,                                 --   clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,  -- reset.reset_n
			address    => mm_interconnect_0_systimer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_systimer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_systimer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_systimer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_systimer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                       --   irq.irq
		);

	mm_interconnect_0 : component raytracing_mm_interconnect_0
		port map (
			altpll_c0_clk                                              => altpll_c0_clk,                                             --                                            altpll_c0.clk
			altpll_c1_clk                                              => altpll_c1_clk,                                             --                                            altpll_c1.clk
			altpll_c3_clk                                              => altpll_c3_clk,                                             --                                            altpll_c3.clk
			clk_50_clk_clk                                             => clk_clk,                                                   --                                           clk_50_clk.clk
			altpll_inclk_interface_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                            --   altpll_inclk_interface_reset_reset_bridge_in_reset.reset
			framereader_clock_master_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                        -- framereader_clock_master_reset_reset_bridge_in_reset.reset
			framereader_clock_reset_reset_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                        --  framereader_clock_reset_reset_reset_bridge_in_reset.reset
			mm_raytracing_0_reset_sink_reset_bridge_in_reset_reset     => rst_controller_003_reset_out_reset,                        --     mm_raytracing_0_reset_sink_reset_bridge_in_reset.reset
			nios2_reset_reset_bridge_in_reset_reset                    => rst_controller_004_reset_out_reset,                        --                    nios2_reset_reset_bridge_in_reset.reset
			framereader_avalon_master_address                          => framereader_avalon_master_address,                         --                            framereader_avalon_master.address
			framereader_avalon_master_waitrequest                      => framereader_avalon_master_waitrequest,                     --                                                     .waitrequest
			framereader_avalon_master_burstcount                       => framereader_avalon_master_burstcount,                      --                                                     .burstcount
			framereader_avalon_master_read                             => framereader_avalon_master_read,                            --                                                     .read
			framereader_avalon_master_readdata                         => framereader_avalon_master_readdata,                        --                                                     .readdata
			framereader_avalon_master_readdatavalid                    => framereader_avalon_master_readdatavalid,                   --                                                     .readdatavalid
			mm_raytracing_0_mm_sdram_master_address                    => mm_raytracing_0_mm_sdram_master_address,                   --                      mm_raytracing_0_mm_sdram_master.address
			mm_raytracing_0_mm_sdram_master_waitrequest                => mm_raytracing_0_mm_sdram_master_waitrequest,               --                                                     .waitrequest
			mm_raytracing_0_mm_sdram_master_write                      => mm_raytracing_0_mm_sdram_master_write,                     --                                                     .write
			mm_raytracing_0_mm_sdram_master_writedata                  => mm_raytracing_0_mm_sdram_master_writedata,                 --                                                     .writedata
			nios2_data_master_address                                  => nios2_data_master_address,                                 --                                    nios2_data_master.address
			nios2_data_master_waitrequest                              => nios2_data_master_waitrequest,                             --                                                     .waitrequest
			nios2_data_master_byteenable                               => nios2_data_master_byteenable,                              --                                                     .byteenable
			nios2_data_master_read                                     => nios2_data_master_read,                                    --                                                     .read
			nios2_data_master_readdata                                 => nios2_data_master_readdata,                                --                                                     .readdata
			nios2_data_master_readdatavalid                            => nios2_data_master_readdatavalid,                           --                                                     .readdatavalid
			nios2_data_master_write                                    => nios2_data_master_write,                                   --                                                     .write
			nios2_data_master_writedata                                => nios2_data_master_writedata,                               --                                                     .writedata
			nios2_data_master_debugaccess                              => nios2_data_master_debugaccess,                             --                                                     .debugaccess
			nios2_instruction_master_address                           => nios2_instruction_master_address,                          --                             nios2_instruction_master.address
			nios2_instruction_master_waitrequest                       => nios2_instruction_master_waitrequest,                      --                                                     .waitrequest
			nios2_instruction_master_read                              => nios2_instruction_master_read,                             --                                                     .read
			nios2_instruction_master_readdata                          => nios2_instruction_master_readdata,                         --                                                     .readdata
			nios2_instruction_master_readdatavalid                     => nios2_instruction_master_readdatavalid,                    --                                                     .readdatavalid
			altpll_pll_slave_address                                   => mm_interconnect_0_altpll_pll_slave_address,                --                                     altpll_pll_slave.address
			altpll_pll_slave_write                                     => mm_interconnect_0_altpll_pll_slave_write,                  --                                                     .write
			altpll_pll_slave_read                                      => mm_interconnect_0_altpll_pll_slave_read,                   --                                                     .read
			altpll_pll_slave_readdata                                  => mm_interconnect_0_altpll_pll_slave_readdata,               --                                                     .readdata
			altpll_pll_slave_writedata                                 => mm_interconnect_0_altpll_pll_slave_writedata,              --                                                     .writedata
			framereader_avalon_slave_address                           => mm_interconnect_0_framereader_avalon_slave_address,        --                             framereader_avalon_slave.address
			framereader_avalon_slave_write                             => mm_interconnect_0_framereader_avalon_slave_write,          --                                                     .write
			framereader_avalon_slave_read                              => mm_interconnect_0_framereader_avalon_slave_read,           --                                                     .read
			framereader_avalon_slave_readdata                          => mm_interconnect_0_framereader_avalon_slave_readdata,       --                                                     .readdata
			framereader_avalon_slave_writedata                         => mm_interconnect_0_framereader_avalon_slave_writedata,      --                                                     .writedata
			jtag_uart_avalon_jtag_slave_address                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                          jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                     .write
			jtag_uart_avalon_jtag_slave_read                           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                     .read
			jtag_uart_avalon_jtag_slave_readdata                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                     .readdata
			jtag_uart_avalon_jtag_slave_writedata                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                     .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                     .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                                     .chipselect
			mm_raytracing_0_mm_nios_slave_address                      => mm_interconnect_0_mm_raytracing_0_mm_nios_slave_address,   --                        mm_raytracing_0_mm_nios_slave.address
			mm_raytracing_0_mm_nios_slave_write                        => mm_interconnect_0_mm_raytracing_0_mm_nios_slave_write,     --                                                     .write
			mm_raytracing_0_mm_nios_slave_writedata                    => mm_interconnect_0_mm_raytracing_0_mm_nios_slave_writedata, --                                                     .writedata
			nios2_debug_mem_slave_address                              => mm_interconnect_0_nios2_debug_mem_slave_address,           --                                nios2_debug_mem_slave.address
			nios2_debug_mem_slave_write                                => mm_interconnect_0_nios2_debug_mem_slave_write,             --                                                     .write
			nios2_debug_mem_slave_read                                 => mm_interconnect_0_nios2_debug_mem_slave_read,              --                                                     .read
			nios2_debug_mem_slave_readdata                             => mm_interconnect_0_nios2_debug_mem_slave_readdata,          --                                                     .readdata
			nios2_debug_mem_slave_writedata                            => mm_interconnect_0_nios2_debug_mem_slave_writedata,         --                                                     .writedata
			nios2_debug_mem_slave_byteenable                           => mm_interconnect_0_nios2_debug_mem_slave_byteenable,        --                                                     .byteenable
			nios2_debug_mem_slave_waitrequest                          => mm_interconnect_0_nios2_debug_mem_slave_waitrequest,       --                                                     .waitrequest
			nios2_debug_mem_slave_debugaccess                          => mm_interconnect_0_nios2_debug_mem_slave_debugaccess,       --                                                     .debugaccess
			onchip_ram_s1_address                                      => mm_interconnect_0_onchip_ram_s1_address,                   --                                        onchip_ram_s1.address
			onchip_ram_s1_write                                        => mm_interconnect_0_onchip_ram_s1_write,                     --                                                     .write
			onchip_ram_s1_readdata                                     => mm_interconnect_0_onchip_ram_s1_readdata,                  --                                                     .readdata
			onchip_ram_s1_writedata                                    => mm_interconnect_0_onchip_ram_s1_writedata,                 --                                                     .writedata
			onchip_ram_s1_byteenable                                   => mm_interconnect_0_onchip_ram_s1_byteenable,                --                                                     .byteenable
			onchip_ram_s1_chipselect                                   => mm_interconnect_0_onchip_ram_s1_chipselect,                --                                                     .chipselect
			onchip_ram_s1_clken                                        => mm_interconnect_0_onchip_ram_s1_clken,                     --                                                     .clken
			sdram_s1_address                                           => mm_interconnect_0_sdram_s1_address,                        --                                             sdram_s1.address
			sdram_s1_write                                             => mm_interconnect_0_sdram_s1_write,                          --                                                     .write
			sdram_s1_read                                              => mm_interconnect_0_sdram_s1_read,                           --                                                     .read
			sdram_s1_readdata                                          => mm_interconnect_0_sdram_s1_readdata,                       --                                                     .readdata
			sdram_s1_writedata                                         => mm_interconnect_0_sdram_s1_writedata,                      --                                                     .writedata
			sdram_s1_byteenable                                        => mm_interconnect_0_sdram_s1_byteenable,                     --                                                     .byteenable
			sdram_s1_readdatavalid                                     => mm_interconnect_0_sdram_s1_readdatavalid,                  --                                                     .readdatavalid
			sdram_s1_waitrequest                                       => mm_interconnect_0_sdram_s1_waitrequest,                    --                                                     .waitrequest
			sdram_s1_chipselect                                        => mm_interconnect_0_sdram_s1_chipselect,                     --                                                     .chipselect
			systimer_s1_address                                        => mm_interconnect_0_systimer_s1_address,                     --                                          systimer_s1.address
			systimer_s1_write                                          => mm_interconnect_0_systimer_s1_write,                       --                                                     .write
			systimer_s1_readdata                                       => mm_interconnect_0_systimer_s1_readdata,                    --                                                     .readdata
			systimer_s1_writedata                                      => mm_interconnect_0_systimer_s1_writedata,                   --                                                     .writedata
			systimer_s1_chipselect                                     => mm_interconnect_0_systimer_s1_chipselect                   --                                                     .chipselect
		);

	irq_mapper : component raytracing_irq_mapper
		port map (
			clk           => altpll_c0_clk,                      --       clk.clk
			reset         => rst_controller_004_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			sender_irq    => nios2_irq_irq                       --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_c1_clk,                      --       receiver_clk.clk
			sender_clk     => altpll_c0_clk,                      --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_004_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	rst_controller : component raytracing_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component raytracing_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_c1_clk,                      --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component raytracing_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => altpll_c0_clk,                          --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component raytracing_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_c3_clk,                      --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component raytracing_rst_controller_004
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,        -- reset_in1.reset
			clk            => altpll_c0_clk,                          --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_004_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_systimer_s1_write_ports_inv <= not mm_interconnect_0_systimer_s1_write;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	ltm_clk_clk <= altpll_c1_clk;

end architecture rtl; -- of raytracing
